`ifndef SER_REF_MODEL_PKG
`define SER_REF_MODEL_PKG

package ser_ref_model_pkg;
    import uvm_pkg::*;
   `include "uvm_macros.svh"
   
   import ser_agent_pkg::*;
   
   `include "ser_ref_model.sv"
   
endpackage

`endif
