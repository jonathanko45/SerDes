`ifndef SER_REF_MODEL
`define SER_REF_MODEL

class ser_ref_model extends uvm_component;
   
    `uvm_component_utils(ser_ref_model);
    
    uvm_analysis_export#(ser_transaction) rm_export;
    uvm_analysis_port#(ser_transaction) rm2sb_port;
    ser_transaction exp_trans, rm_trans;
    uvm_tlm_analysis_fifo#(ser_transaction) rm_exp_fifo;
    uvm_queue#(int) rm_queue = uvm_queue_pool::get_global("queue_key_rm");
    int RD;
    
    function new(string name = "ser_ref_model", uvm_component parent);
        super.new(name, parent);
    endfunction: new
    
    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        rm_export = new("rm_export", this);
        rm2sb_port = new("rm2sb_port", this);
        rm_exp_fifo = new("rm_exp_fifo", this);
        if(!uvm_config_db#(int)::get(this, "", "running_disparity", RD))
            `uvm_fatal("NO RD", {"Running Disparity must be set for: ", get_full_name(), ".RD"})
    endfunction: build_phase
    
    function void connect_phase(uvm_phase phase);
        super.connect_phase(phase);
        rm_export.connect(rm_exp_fifo.analysis_export);
    endfunction: connect_phase
    
    task run_phase(uvm_phase phase);
        forever begin
            rm_exp_fifo.get(rm_trans);
            get_expected_transaction(rm_trans);
        end
     endtask
     
     task get_expected_transaction(ser_transaction rm_trans);
        this.exp_trans = rm_trans;
        exp_trans.in_RD = RD;
        if (RD == 2'sb11) begin
            case (exp_trans.in_data)
                8'b00000000 : exp_trans.out_10b = 10'b1001110100;
                8'b00000001 : exp_trans.out_10b = 10'b0111010100;
                8'b00000010 : exp_trans.out_10b = 10'b1011010100;
                8'b00000011 : exp_trans.out_10b = 10'b1100011011;
                8'b00000100 : exp_trans.out_10b = 10'b1101010100;
                8'b00000101 : exp_trans.out_10b = 10'b1010011011;
                8'b00000110 : exp_trans.out_10b = 10'b0110011011;
                8'b00000111 : exp_trans.out_10b = 10'b1110001011;
                8'b00001000 : exp_trans.out_10b = 10'b1110010100;
                8'b00001001 : exp_trans.out_10b = 10'b1001011011;
                8'b00001010 : exp_trans.out_10b = 10'b0101011011;
                8'b00001011 : exp_trans.out_10b = 10'b1101001011;
                8'b00001100 : exp_trans.out_10b = 10'b0011011011;
                8'b00001101 : exp_trans.out_10b = 10'b1011001011;
                8'b00001110 : exp_trans.out_10b = 10'b0111001011;
                8'b00001111 : exp_trans.out_10b = 10'b0101110100;
                8'b00010000 : exp_trans.out_10b = 10'b0110110100;
                8'b00010001 : exp_trans.out_10b = 10'b1000111011;
                8'b00010010 : exp_trans.out_10b = 10'b0100111011;
                8'b00010011 : exp_trans.out_10b = 10'b1100101011;
                8'b00010100 : exp_trans.out_10b = 10'b0010111011;
                8'b00010101 : exp_trans.out_10b = 10'b1010101011;
                8'b00010110 : exp_trans.out_10b = 10'b0110101011;
                8'b00010111 : exp_trans.out_10b = 10'b1110100100;
                8'b00011000 : exp_trans.out_10b = 10'b1100110100;
                8'b00011001 : exp_trans.out_10b = 10'b1001101011;
                8'b00011010 : exp_trans.out_10b = 10'b0101101011;
                8'b00011011 : exp_trans.out_10b = 10'b1101100100;
                8'b00011100 : exp_trans.out_10b = 10'b0011101011;
                8'b00011101 : exp_trans.out_10b = 10'b1011100100;
                8'b00011110 : exp_trans.out_10b = 10'b0111100100;
                8'b00011111 : exp_trans.out_10b = 10'b1010110100;
                8'b00100000 : exp_trans.out_10b = 10'b1001111001;
                8'b00100001 : exp_trans.out_10b = 10'b0111011001;
                8'b00100010 : exp_trans.out_10b = 10'b1011011001;
                8'b00100011 : exp_trans.out_10b = 10'b1100011001;
                8'b00100100 : exp_trans.out_10b = 10'b1101011001;
                8'b00100101 : exp_trans.out_10b = 10'b1010011001;
                8'b00100110 : exp_trans.out_10b = 10'b0110011001;
                8'b00100111 : exp_trans.out_10b = 10'b1110001001;
                8'b00101000 : exp_trans.out_10b = 10'b1110011001;
                8'b00101001 : exp_trans.out_10b = 10'b1001011001;
                8'b00101010 : exp_trans.out_10b = 10'b0101011001;
                8'b00101011 : exp_trans.out_10b = 10'b1101001001;
                8'b00101100 : exp_trans.out_10b = 10'b0011011001;
                8'b00101101 : exp_trans.out_10b = 10'b1011001001;
                8'b00101110 : exp_trans.out_10b = 10'b0111001001;
                8'b00101111 : exp_trans.out_10b = 10'b0101111001;
                8'b00110000 : exp_trans.out_10b = 10'b0110111001;
                8'b00110001 : exp_trans.out_10b = 10'b1000111001;
                8'b00110010 : exp_trans.out_10b = 10'b0100111001;
                8'b00110011 : exp_trans.out_10b = 10'b1100101001;
                8'b00110100 : exp_trans.out_10b = 10'b0010111001;
                8'b00110101 : exp_trans.out_10b = 10'b1010101001;
                8'b00110110 : exp_trans.out_10b = 10'b0110101001;
                8'b00110111 : exp_trans.out_10b = 10'b1110101001;
                8'b00111000 : exp_trans.out_10b = 10'b1100111001;
                8'b00111001 : exp_trans.out_10b = 10'b1001101001;
                8'b00111010 : exp_trans.out_10b = 10'b0101101001;
                8'b00111011 : exp_trans.out_10b = 10'b1101101001;
                8'b00111100 : exp_trans.out_10b = 10'b0011101001;
                8'b00111101 : exp_trans.out_10b = 10'b1011101001;
                8'b00111110 : exp_trans.out_10b = 10'b0111101001;
                8'b00111111 : exp_trans.out_10b = 10'b1010111001;
                8'b01000000 : exp_trans.out_10b = 10'b1001110101;
                8'b01000001 : exp_trans.out_10b = 10'b0111010101;
                8'b01000010 : exp_trans.out_10b = 10'b1011010101;
                8'b01000011 : exp_trans.out_10b = 10'b1100010101;
                8'b01000100 : exp_trans.out_10b = 10'b1101010101;
                8'b01000101 : exp_trans.out_10b = 10'b1010010101;
                8'b01000110 : exp_trans.out_10b = 10'b0110010101;
                8'b01000111 : exp_trans.out_10b = 10'b1110000101;
                8'b01001000 : exp_trans.out_10b = 10'b1110010101;
                8'b01001001 : exp_trans.out_10b = 10'b1001010101;
                8'b01001010 : exp_trans.out_10b = 10'b0101010101;
                8'b01001011 : exp_trans.out_10b = 10'b1101000101;
                8'b01001100 : exp_trans.out_10b = 10'b0011010101;
                8'b01001101 : exp_trans.out_10b = 10'b1011000101;
                8'b01001110 : exp_trans.out_10b = 10'b0111000101;
                8'b01001111 : exp_trans.out_10b = 10'b0101110101;
                8'b01010000 : exp_trans.out_10b = 10'b0110110101;
                8'b01010001 : exp_trans.out_10b = 10'b1000110101;
                8'b01010010 : exp_trans.out_10b = 10'b0100110101;
                8'b01010011 : exp_trans.out_10b = 10'b1100100101;
                8'b01010100 : exp_trans.out_10b = 10'b0010110101;
                8'b01010101 : exp_trans.out_10b = 10'b1010100101;
                8'b01010110 : exp_trans.out_10b = 10'b0110100101;
                8'b01010111 : exp_trans.out_10b = 10'b1110100101;
                8'b01011000 : exp_trans.out_10b = 10'b1100110101;
                8'b01011001 : exp_trans.out_10b = 10'b1001100101;
                8'b01011010 : exp_trans.out_10b = 10'b0101100101;
                8'b01011011 : exp_trans.out_10b = 10'b1101100101;
                8'b01011100 : exp_trans.out_10b = 10'b0011100101;
                8'b01011101 : exp_trans.out_10b = 10'b1011100101;
                8'b01011110 : exp_trans.out_10b = 10'b0111100101;
                8'b01011111 : exp_trans.out_10b = 10'b1010110101;
                8'b01100000 : exp_trans.out_10b = 10'b1001110011;
                8'b01100001 : exp_trans.out_10b = 10'b0111010011;
                8'b01100010 : exp_trans.out_10b = 10'b1011010011;
                8'b01100011 : exp_trans.out_10b = 10'b1100011100;
                8'b01100100 : exp_trans.out_10b = 10'b1101010011;
                8'b01100101 : exp_trans.out_10b = 10'b1010011100;
                8'b01100110 : exp_trans.out_10b = 10'b0110011100;
                8'b01100111 : exp_trans.out_10b = 10'b1110001100;
                8'b01101000 : exp_trans.out_10b = 10'b1110010011;
                8'b01101001 : exp_trans.out_10b = 10'b1001011100;
                8'b01101010 : exp_trans.out_10b = 10'b0101011100;
                8'b01101011 : exp_trans.out_10b = 10'b1101001100;
                8'b01101100 : exp_trans.out_10b = 10'b0011011100;
                8'b01101101 : exp_trans.out_10b = 10'b1011001100;
                8'b01101110 : exp_trans.out_10b = 10'b0111001100;
                8'b01101111 : exp_trans.out_10b = 10'b0101110011;
                8'b01110000 : exp_trans.out_10b = 10'b0110110011;
                8'b01110001 : exp_trans.out_10b = 10'b1000111100;
                8'b01110010 : exp_trans.out_10b = 10'b0100111100;
                8'b01110011 : exp_trans.out_10b = 10'b1100101100;
                8'b01110100 : exp_trans.out_10b = 10'b0010111100;
                8'b01110101 : exp_trans.out_10b = 10'b1010101100;
                8'b01110110 : exp_trans.out_10b = 10'b0110101100;
                8'b01110111 : exp_trans.out_10b = 10'b1110100011;
                8'b01111000 : exp_trans.out_10b = 10'b1100110011;
                8'b01111001 : exp_trans.out_10b = 10'b1001101100;
                8'b01111010 : exp_trans.out_10b = 10'b0101101100;
                8'b01111011 : exp_trans.out_10b = 10'b1101100011;
                8'b01111100 : exp_trans.out_10b = 10'b0011101100;
                8'b01111101 : exp_trans.out_10b = 10'b1011100011;
                8'b01111110 : exp_trans.out_10b = 10'b0111100011;
                8'b01111111 : exp_trans.out_10b = 10'b1010110011;
                8'b10000000 : exp_trans.out_10b = 10'b1001110010;
                8'b10000001 : exp_trans.out_10b = 10'b0111010010;
                8'b10000010 : exp_trans.out_10b = 10'b1011010010;
                8'b10000011 : exp_trans.out_10b = 10'b1100011101;
                8'b10000100 : exp_trans.out_10b = 10'b1101010010;
                8'b10000101 : exp_trans.out_10b = 10'b1010011101;
                8'b10000110 : exp_trans.out_10b = 10'b0110011101;
                8'b10000111 : exp_trans.out_10b = 10'b1110001101;
                8'b10001000 : exp_trans.out_10b = 10'b1110010010;
                8'b10001001 : exp_trans.out_10b = 10'b1001011101;
                8'b10001010 : exp_trans.out_10b = 10'b0101011101;
                8'b10001011 : exp_trans.out_10b = 10'b1101001101;
                8'b10001100 : exp_trans.out_10b = 10'b0011011101;
                8'b10001101 : exp_trans.out_10b = 10'b1011001101;
                8'b10001110 : exp_trans.out_10b = 10'b0111001101;
                8'b10001111 : exp_trans.out_10b = 10'b0101110010;
                8'b10010000 : exp_trans.out_10b = 10'b0110110010;
                8'b10010001 : exp_trans.out_10b = 10'b1000111101;
                8'b10010010 : exp_trans.out_10b = 10'b0100111101;
                8'b10010011 : exp_trans.out_10b = 10'b1100101101;
                8'b10010100 : exp_trans.out_10b = 10'b0010111101;
                8'b10010101 : exp_trans.out_10b = 10'b1010101101;
                8'b10010110 : exp_trans.out_10b = 10'b0110101101;
                8'b10010111 : exp_trans.out_10b = 10'b1110100010;
                8'b10011000 : exp_trans.out_10b = 10'b1100110010;
                8'b10011001 : exp_trans.out_10b = 10'b1001101101;
                8'b10011010 : exp_trans.out_10b = 10'b0101101101;
                8'b10011011 : exp_trans.out_10b = 10'b1101100010;
                8'b10011100 : exp_trans.out_10b = 10'b0011101101;
                8'b10011101 : exp_trans.out_10b = 10'b1011100010;
                8'b10011110 : exp_trans.out_10b = 10'b0111100010;
                8'b10011111 : exp_trans.out_10b = 10'b1010110010;
                8'b10100000 : exp_trans.out_10b = 10'b1001111010;
                8'b10100001 : exp_trans.out_10b = 10'b0111011010;
                8'b10100010 : exp_trans.out_10b = 10'b1011011010;
                8'b10100011 : exp_trans.out_10b = 10'b1100011010;
                8'b10100100 : exp_trans.out_10b = 10'b1101011010;
                8'b10100101 : exp_trans.out_10b = 10'b1010011010;
                8'b10100110 : exp_trans.out_10b = 10'b0110011010;
                8'b10100111 : exp_trans.out_10b = 10'b1110001010;
                8'b10101000 : exp_trans.out_10b = 10'b1110011010;
                8'b10101001 : exp_trans.out_10b = 10'b1001011010;
                8'b10101010 : exp_trans.out_10b = 10'b0101011010;
                8'b10101011 : exp_trans.out_10b = 10'b1101001010;
                8'b10101100 : exp_trans.out_10b = 10'b0011011010;
                8'b10101101 : exp_trans.out_10b = 10'b1011001010;
                8'b10101110 : exp_trans.out_10b = 10'b0111001010;
                8'b10101111 : exp_trans.out_10b = 10'b0101111010;
                8'b10110000 : exp_trans.out_10b = 10'b0110111010;
                8'b10110001 : exp_trans.out_10b = 10'b1000111010;
                8'b10110010 : exp_trans.out_10b = 10'b0100111010;
                8'b10110011 : exp_trans.out_10b = 10'b1100101010;
                8'b10110100 : exp_trans.out_10b = 10'b0010111010;
                8'b10110101 : exp_trans.out_10b = 10'b1010101010;
                8'b10110110 : exp_trans.out_10b = 10'b0110101010;
                8'b10110111 : exp_trans.out_10b = 10'b1110101010;
                8'b10111000 : exp_trans.out_10b = 10'b1100111010;
                8'b10111001 : exp_trans.out_10b = 10'b1001101010;
                8'b10111010 : exp_trans.out_10b = 10'b0101101010;
                8'b10111011 : exp_trans.out_10b = 10'b1101101010;
                8'b10111100 : exp_trans.out_10b = 10'b0011101010;
                8'b10111101 : exp_trans.out_10b = 10'b1011101010;
                8'b10111110 : exp_trans.out_10b = 10'b0111101010;
                8'b10111111 : exp_trans.out_10b = 10'b1010111010;
                8'b11000000 : exp_trans.out_10b = 10'b1001110110;
                8'b11000001 : exp_trans.out_10b = 10'b0111010110;
                8'b11000010 : exp_trans.out_10b = 10'b1011010110;
                8'b11000011 : exp_trans.out_10b = 10'b1100010110;
                8'b11000100 : exp_trans.out_10b = 10'b1101010110;
                8'b11000101 : exp_trans.out_10b = 10'b1010010110;
                8'b11000110 : exp_trans.out_10b = 10'b0110010110;
                8'b11000111 : exp_trans.out_10b = 10'b1110000110;
                8'b11001000 : exp_trans.out_10b = 10'b1110010110;
                8'b11001001 : exp_trans.out_10b = 10'b1001010110;
                8'b11001010 : exp_trans.out_10b = 10'b0101010110;
                8'b11001011 : exp_trans.out_10b = 10'b1101000110;
                8'b11001100 : exp_trans.out_10b = 10'b0011010110;
                8'b11001101 : exp_trans.out_10b = 10'b1011000110;
                8'b11001110 : exp_trans.out_10b = 10'b0111000110;
                8'b11001111 : exp_trans.out_10b = 10'b0101110110;
                8'b11010000 : exp_trans.out_10b = 10'b0110110110;
                8'b11010001 : exp_trans.out_10b = 10'b1000110110;
                8'b11010010 : exp_trans.out_10b = 10'b0100110110;
                8'b11010011 : exp_trans.out_10b = 10'b1100100110;
                8'b11010100 : exp_trans.out_10b = 10'b0010110110;
                8'b11010101 : exp_trans.out_10b = 10'b1010100110;
                8'b11010110 : exp_trans.out_10b = 10'b0110100110;
                8'b11010111 : exp_trans.out_10b = 10'b1110100110;
                8'b11011000 : exp_trans.out_10b = 10'b1100110110;
                8'b11011001 : exp_trans.out_10b = 10'b1001100110;
                8'b11011010 : exp_trans.out_10b = 10'b0101100110;
                8'b11011011 : exp_trans.out_10b = 10'b1101100110;
                8'b11011100 : exp_trans.out_10b = 10'b0011100110;
                8'b11011101 : exp_trans.out_10b = 10'b1011100110;
                8'b11011110 : exp_trans.out_10b = 10'b0111100110;
                8'b11011111 : exp_trans.out_10b = 10'b1010110110;
                8'b11100000 : exp_trans.out_10b = 10'b1001110001;
                8'b11100001 : exp_trans.out_10b = 10'b0111010001;
                8'b11100010 : exp_trans.out_10b = 10'b1011010001;
                8'b11100011 : exp_trans.out_10b = 10'b1100011110;
                8'b11100100 : exp_trans.out_10b = 10'b1101010001;
                8'b11100101 : exp_trans.out_10b = 10'b1010011110;
                8'b11100110 : exp_trans.out_10b = 10'b0110011110;
                8'b11100111 : exp_trans.out_10b = 10'b1110001110;
                8'b11101000 : exp_trans.out_10b = 10'b1110010001;
                8'b11101001 : exp_trans.out_10b = 10'b1001011110;
                8'b11101010 : exp_trans.out_10b = 10'b0101011110;
                8'b11101011 : exp_trans.out_10b = 10'b1101001110;
                8'b11101100 : exp_trans.out_10b = 10'b0011011110;
                8'b11101101 : exp_trans.out_10b = 10'b1011001110;
                8'b11101110 : exp_trans.out_10b = 10'b0111001110;
                8'b11101111 : exp_trans.out_10b = 10'b0101110001;
                8'b11110000 : exp_trans.out_10b = 10'b0110110001;
                8'b11110001 : exp_trans.out_10b = 10'b1000110111;
                8'b11110010 : exp_trans.out_10b = 10'b0100110111;
                8'b11110011 : exp_trans.out_10b = 10'b1100101110;
                8'b11110100 : exp_trans.out_10b = 10'b0010110111;
                8'b11110101 : exp_trans.out_10b = 10'b1010101110;
                8'b11110110 : exp_trans.out_10b = 10'b0110101110;
                8'b11110111 : exp_trans.out_10b = 10'b1110100001;
                8'b11111000 : exp_trans.out_10b = 10'b1100110001;
                8'b11111001 : exp_trans.out_10b = 10'b1001101110;
                8'b11111010 : exp_trans.out_10b = 10'b0101101110;
                8'b11111011 : exp_trans.out_10b = 10'b1101100001;
                8'b11111100 : exp_trans.out_10b = 10'b0011101110;
                8'b11111101 : exp_trans.out_10b = 10'b1011100001;
                8'b11111110 : exp_trans.out_10b = 10'b0111100001;
                8'b11111111 : exp_trans.out_10b = 10'b1010110001;
                default : exp_trans.out_10b = 10'b0000000000;
            endcase
        end else if(RD == 2'sb01) begin
            case (exp_trans.in_data)
                8'b00000000 : exp_trans.out_10b = 10'b0110001011;
                8'b00000001 : exp_trans.out_10b = 10'b1000101011;
                8'b00000010 : exp_trans.out_10b = 10'b0100101011;
                8'b00000011 : exp_trans.out_10b = 10'b1100010100;
                8'b00000100 : exp_trans.out_10b = 10'b0010101011;
                8'b00000101 : exp_trans.out_10b = 10'b1010010100;
                8'b00000110 : exp_trans.out_10b = 10'b0110010100;
                8'b00000111 : exp_trans.out_10b = 10'b0001110100;
                8'b00001000 : exp_trans.out_10b = 10'b0001101011;
                8'b00001001 : exp_trans.out_10b = 10'b1001010100;
                8'b00001010 : exp_trans.out_10b = 10'b0101010100;
                8'b00001011 : exp_trans.out_10b = 10'b1101000100;
                8'b00001100 : exp_trans.out_10b = 10'b0011010100;
                8'b00001101 : exp_trans.out_10b = 10'b1011000100;
                8'b00001110 : exp_trans.out_10b = 10'b0111000100;
                8'b00001111 : exp_trans.out_10b = 10'b1010001011;
                8'b00010000 : exp_trans.out_10b = 10'b1001001011;
                8'b00010001 : exp_trans.out_10b = 10'b1000110100;
                8'b00010010 : exp_trans.out_10b = 10'b0100110100;
                8'b00010011 : exp_trans.out_10b = 10'b1100100100;
                8'b00010100 : exp_trans.out_10b = 10'b0010110100;
                8'b00010101 : exp_trans.out_10b = 10'b1010100100;
                8'b00010110 : exp_trans.out_10b = 10'b0110100100;
                8'b00010111 : exp_trans.out_10b = 10'b0001011011;
                8'b00011000 : exp_trans.out_10b = 10'b0011001011;
                8'b00011001 : exp_trans.out_10b = 10'b1001100100;
                8'b00011010 : exp_trans.out_10b = 10'b0101100100;
                8'b00011011 : exp_trans.out_10b = 10'b0010011011;
                8'b00011100 : exp_trans.out_10b = 10'b0011100100;
                8'b00011101 : exp_trans.out_10b = 10'b0100011011;
                8'b00011110 : exp_trans.out_10b = 10'b1000011011;
                8'b00011111 : exp_trans.out_10b = 10'b0101001011;
                8'b00100000 : exp_trans.out_10b = 10'b0110001001;
                8'b00100001 : exp_trans.out_10b = 10'b1000101001;
                8'b00100010 : exp_trans.out_10b = 10'b0100101001;
                8'b00100011 : exp_trans.out_10b = 10'b1100011001;
                8'b00100100 : exp_trans.out_10b = 10'b0010101001;
                8'b00100101 : exp_trans.out_10b = 10'b1010011001;
                8'b00100110 : exp_trans.out_10b = 10'b0110011001;
                8'b00100111 : exp_trans.out_10b = 10'b0001111001;
                8'b00101000 : exp_trans.out_10b = 10'b0001101001;
                8'b00101001 : exp_trans.out_10b = 10'b1001011001;
                8'b00101010 : exp_trans.out_10b = 10'b0101011001;
                8'b00101011 : exp_trans.out_10b = 10'b1101001001;
                8'b00101100 : exp_trans.out_10b = 10'b0011011001;
                8'b00101101 : exp_trans.out_10b = 10'b1011001001;
                8'b00101110 : exp_trans.out_10b = 10'b0111001001;
                8'b00101111 : exp_trans.out_10b = 10'b1010001001;
                8'b00110000 : exp_trans.out_10b = 10'b1001001001;
                8'b00110001 : exp_trans.out_10b = 10'b1000111001;
                8'b00110010 : exp_trans.out_10b = 10'b0100111001;
                8'b00110011 : exp_trans.out_10b = 10'b1100101001;
                8'b00110100 : exp_trans.out_10b = 10'b0010111001;
                8'b00110101 : exp_trans.out_10b = 10'b1010101001;
                8'b00110110 : exp_trans.out_10b = 10'b0110101001;
                8'b00110111 : exp_trans.out_10b = 10'b0001011001;
                8'b00111000 : exp_trans.out_10b = 10'b0011001001;
                8'b00111001 : exp_trans.out_10b = 10'b1001101001;
                8'b00111010 : exp_trans.out_10b = 10'b0101101001;
                8'b00111011 : exp_trans.out_10b = 10'b0010011001;
                8'b00111100 : exp_trans.out_10b = 10'b0011101001;
                8'b00111101 : exp_trans.out_10b = 10'b0100011001;
                8'b00111110 : exp_trans.out_10b = 10'b1000011001;
                8'b00111111 : exp_trans.out_10b = 10'b0101001001;
                8'b01000000 : exp_trans.out_10b = 10'b0110000101;
                8'b01000001 : exp_trans.out_10b = 10'b1000100101;
                8'b01000010 : exp_trans.out_10b = 10'b0100100101;
                8'b01000011 : exp_trans.out_10b = 10'b1100010101;
                8'b01000100 : exp_trans.out_10b = 10'b0010100101;
                8'b01000101 : exp_trans.out_10b = 10'b1010010101;
                8'b01000110 : exp_trans.out_10b = 10'b0110010101;
                8'b01000111 : exp_trans.out_10b = 10'b0001110101;
                8'b01001000 : exp_trans.out_10b = 10'b0001100101;
                8'b01001001 : exp_trans.out_10b = 10'b1001010101;
                8'b01001010 : exp_trans.out_10b = 10'b0101010101;
                8'b01001011 : exp_trans.out_10b = 10'b1101000101;
                8'b01001100 : exp_trans.out_10b = 10'b0011010101;
                8'b01001101 : exp_trans.out_10b = 10'b1011000101;
                8'b01001110 : exp_trans.out_10b = 10'b0111000101;
                8'b01001111 : exp_trans.out_10b = 10'b1010000101;
                8'b01010000 : exp_trans.out_10b = 10'b1001000101;
                8'b01010001 : exp_trans.out_10b = 10'b1000110101;
                8'b01010010 : exp_trans.out_10b = 10'b0100110101;
                8'b01010011 : exp_trans.out_10b = 10'b1100100101;
                8'b01010100 : exp_trans.out_10b = 10'b0010110101;
                8'b01010101 : exp_trans.out_10b = 10'b1010100101;
                8'b01010110 : exp_trans.out_10b = 10'b0110100101;
                8'b01010111 : exp_trans.out_10b = 10'b0001010101;
                8'b01011000 : exp_trans.out_10b = 10'b0011000101;
                8'b01011001 : exp_trans.out_10b = 10'b1001100101;
                8'b01011010 : exp_trans.out_10b = 10'b0101100101;
                8'b01011011 : exp_trans.out_10b = 10'b0010010101;
                8'b01011100 : exp_trans.out_10b = 10'b0011100101;
                8'b01011101 : exp_trans.out_10b = 10'b0100010101;
                8'b01011110 : exp_trans.out_10b = 10'b1000010101;
                8'b01011111 : exp_trans.out_10b = 10'b0101000101;
                8'b01100000 : exp_trans.out_10b = 10'b0110001100;
                8'b01100001 : exp_trans.out_10b = 10'b1000101100;
                8'b01100010 : exp_trans.out_10b = 10'b0100101100;
                8'b01100011 : exp_trans.out_10b = 10'b1100010011;
                8'b01100100 : exp_trans.out_10b = 10'b0010101100;
                8'b01100101 : exp_trans.out_10b = 10'b1010010011;
                8'b01100110 : exp_trans.out_10b = 10'b0110010011;
                8'b01100111 : exp_trans.out_10b = 10'b0001110011;
                8'b01101000 : exp_trans.out_10b = 10'b0001101100;
                8'b01101001 : exp_trans.out_10b = 10'b1001010011;
                8'b01101010 : exp_trans.out_10b = 10'b0101010011;
                8'b01101011 : exp_trans.out_10b = 10'b1101000011;
                8'b01101100 : exp_trans.out_10b = 10'b0011010011;
                8'b01101101 : exp_trans.out_10b = 10'b1011000011;
                8'b01101110 : exp_trans.out_10b = 10'b0111000011;
                8'b01101111 : exp_trans.out_10b = 10'b1010001100;
                8'b01110000 : exp_trans.out_10b = 10'b1001001100;
                8'b01110001 : exp_trans.out_10b = 10'b1000110011;
                8'b01110010 : exp_trans.out_10b = 10'b0100110011;
                8'b01110011 : exp_trans.out_10b = 10'b1100100011;
                8'b01110100 : exp_trans.out_10b = 10'b0010110011;
                8'b01110101 : exp_trans.out_10b = 10'b1010100011;
                8'b01110110 : exp_trans.out_10b = 10'b0110100011;
                8'b01110111 : exp_trans.out_10b = 10'b0001011100;
                8'b01111000 : exp_trans.out_10b = 10'b0011001100;
                8'b01111001 : exp_trans.out_10b = 10'b1001100011;
                8'b01111010 : exp_trans.out_10b = 10'b0101100011;
                8'b01111011 : exp_trans.out_10b = 10'b0010011100;
                8'b01111100 : exp_trans.out_10b = 10'b0011100011;
                8'b01111101 : exp_trans.out_10b = 10'b0100011100;
                8'b01111110 : exp_trans.out_10b = 10'b1000011100;
                8'b01111111 : exp_trans.out_10b = 10'b0101001100;
                8'b10000000 : exp_trans.out_10b = 10'b0110001101;
                8'b10000001 : exp_trans.out_10b = 10'b1000101101;
                8'b10000010 : exp_trans.out_10b = 10'b0100101101;
                8'b10000011 : exp_trans.out_10b = 10'b1100010010;
                8'b10000100 : exp_trans.out_10b = 10'b0010101101;
                8'b10000101 : exp_trans.out_10b = 10'b1010010010;
                8'b10000110 : exp_trans.out_10b = 10'b0110010010;
                8'b10000111 : exp_trans.out_10b = 10'b0001110010;
                8'b10001000 : exp_trans.out_10b = 10'b0001101101;
                8'b10001001 : exp_trans.out_10b = 10'b1001010010;
                8'b10001010 : exp_trans.out_10b = 10'b0101010010;
                8'b10001011 : exp_trans.out_10b = 10'b1101000010;
                8'b10001100 : exp_trans.out_10b = 10'b0011010010;
                8'b10001101 : exp_trans.out_10b = 10'b1011000010;
                8'b10001110 : exp_trans.out_10b = 10'b0111000010;
                8'b10001111 : exp_trans.out_10b = 10'b1010001101;
                8'b10010000 : exp_trans.out_10b = 10'b1001001101;
                8'b10010001 : exp_trans.out_10b = 10'b1000110010;
                8'b10010010 : exp_trans.out_10b = 10'b0100110010;
                8'b10010011 : exp_trans.out_10b = 10'b1100100010;
                8'b10010100 : exp_trans.out_10b = 10'b0010110010;
                8'b10010101 : exp_trans.out_10b = 10'b1010100010;
                8'b10010110 : exp_trans.out_10b = 10'b0110100010;
                8'b10010111 : exp_trans.out_10b = 10'b0001011101;
                8'b10011000 : exp_trans.out_10b = 10'b0011001101;
                8'b10011001 : exp_trans.out_10b = 10'b1001100010;
                8'b10011010 : exp_trans.out_10b = 10'b0101100010;
                8'b10011011 : exp_trans.out_10b = 10'b0010011101;
                8'b10011100 : exp_trans.out_10b = 10'b0011100010;
                8'b10011101 : exp_trans.out_10b = 10'b0100011101;
                8'b10011110 : exp_trans.out_10b = 10'b1000011101;
                8'b10011111 : exp_trans.out_10b = 10'b0101001101;
                8'b10100000 : exp_trans.out_10b = 10'b0110001010;
                8'b10100001 : exp_trans.out_10b = 10'b1000101010;
                8'b10100010 : exp_trans.out_10b = 10'b0100101010;
                8'b10100011 : exp_trans.out_10b = 10'b1100011010;
                8'b10100100 : exp_trans.out_10b = 10'b0010101010;
                8'b10100101 : exp_trans.out_10b = 10'b1010011010;
                8'b10100110 : exp_trans.out_10b = 10'b0110011010;
                8'b10100111 : exp_trans.out_10b = 10'b0001111010;
                8'b10101000 : exp_trans.out_10b = 10'b0001101010;
                8'b10101001 : exp_trans.out_10b = 10'b1001011010;
                8'b10101010 : exp_trans.out_10b = 10'b0101011010;
                8'b10101011 : exp_trans.out_10b = 10'b1101001010;
                8'b10101100 : exp_trans.out_10b = 10'b0011011010;
                8'b10101101 : exp_trans.out_10b = 10'b1011001010;
                8'b10101110 : exp_trans.out_10b = 10'b0111001010;
                8'b10101111 : exp_trans.out_10b = 10'b1010001010;
                8'b10110000 : exp_trans.out_10b = 10'b1001001010;
                8'b10110001 : exp_trans.out_10b = 10'b1000111010;
                8'b10110010 : exp_trans.out_10b = 10'b0100111010;
                8'b10110011 : exp_trans.out_10b = 10'b1100101010;
                8'b10110100 : exp_trans.out_10b = 10'b0010111010;
                8'b10110101 : exp_trans.out_10b = 10'b1010101010;
                8'b10110110 : exp_trans.out_10b = 10'b0110101010;
                8'b10110111 : exp_trans.out_10b = 10'b0001011010;
                8'b10111000 : exp_trans.out_10b = 10'b0011001010;
                8'b10111001 : exp_trans.out_10b = 10'b1001101010;
                8'b10111010 : exp_trans.out_10b = 10'b0101101010;
                8'b10111011 : exp_trans.out_10b = 10'b0010011010;
                8'b10111100 : exp_trans.out_10b = 10'b0011101010;
                8'b10111101 : exp_trans.out_10b = 10'b0100011010;
                8'b10111110 : exp_trans.out_10b = 10'b1000011010;
                8'b10111111 : exp_trans.out_10b = 10'b0101001010;
                8'b11000000 : exp_trans.out_10b = 10'b0110000110;
                8'b11000001 : exp_trans.out_10b = 10'b1000100110;
                8'b11000010 : exp_trans.out_10b = 10'b0100100110;
                8'b11000011 : exp_trans.out_10b = 10'b1100010110;
                8'b11000100 : exp_trans.out_10b = 10'b0010100110;
                8'b11000101 : exp_trans.out_10b = 10'b1010010110;
                8'b11000110 : exp_trans.out_10b = 10'b0110010110;
                8'b11000111 : exp_trans.out_10b = 10'b0001110110;
                8'b11001000 : exp_trans.out_10b = 10'b0001100110;
                8'b11001001 : exp_trans.out_10b = 10'b1001010110;
                8'b11001010 : exp_trans.out_10b = 10'b0101010110;
                8'b11001011 : exp_trans.out_10b = 10'b1101000110;
                8'b11001100 : exp_trans.out_10b = 10'b0011010110;
                8'b11001101 : exp_trans.out_10b = 10'b1011000110;
                8'b11001110 : exp_trans.out_10b = 10'b0111000110;
                8'b11001111 : exp_trans.out_10b = 10'b1010000110;
                8'b11010000 : exp_trans.out_10b = 10'b1001000110;
                8'b11010001 : exp_trans.out_10b = 10'b1000110110;
                8'b11010010 : exp_trans.out_10b = 10'b0100110110;
                8'b11010011 : exp_trans.out_10b = 10'b1100100110;
                8'b11010100 : exp_trans.out_10b = 10'b0010110110;
                8'b11010101 : exp_trans.out_10b = 10'b1010100110;
                8'b11010110 : exp_trans.out_10b = 10'b0110100110;
                8'b11010111 : exp_trans.out_10b = 10'b0001010110;
                8'b11011000 : exp_trans.out_10b = 10'b0011000110;
                8'b11011001 : exp_trans.out_10b = 10'b1001100110;
                8'b11011010 : exp_trans.out_10b = 10'b0101100110;
                8'b11011011 : exp_trans.out_10b = 10'b0010010110;
                8'b11011100 : exp_trans.out_10b = 10'b0011100110;
                8'b11011101 : exp_trans.out_10b = 10'b0100010110;
                8'b11011110 : exp_trans.out_10b = 10'b1000010110;
                8'b11011111 : exp_trans.out_10b = 10'b0101000110;
                8'b11100000 : exp_trans.out_10b = 10'b0110001110;
                8'b11100001 : exp_trans.out_10b = 10'b1000101110;
                8'b11100010 : exp_trans.out_10b = 10'b0100101110;
                8'b11100011 : exp_trans.out_10b = 10'b1100010001;
                8'b11100100 : exp_trans.out_10b = 10'b0010101110;
                8'b11100101 : exp_trans.out_10b = 10'b1010010001;
                8'b11100110 : exp_trans.out_10b = 10'b0110010001;
                8'b11100111 : exp_trans.out_10b = 10'b0001110001;
                8'b11101000 : exp_trans.out_10b = 10'b0001101110;
                8'b11101001 : exp_trans.out_10b = 10'b1001010001;
                8'b11101010 : exp_trans.out_10b = 10'b0101010001;
                8'b11101011 : exp_trans.out_10b = 10'b1101001000;
                8'b11101100 : exp_trans.out_10b = 10'b0011010001;
                8'b11101101 : exp_trans.out_10b = 10'b1011001000;
                8'b11101110 : exp_trans.out_10b = 10'b0111001000;
                8'b11101111 : exp_trans.out_10b = 10'b1010001110;
                8'b11110000 : exp_trans.out_10b = 10'b1001001110;
                8'b11110001 : exp_trans.out_10b = 10'b1000110001;
                8'b11110010 : exp_trans.out_10b = 10'b0100110001;
                8'b11110011 : exp_trans.out_10b = 10'b1100100001;
                8'b11110100 : exp_trans.out_10b = 10'b0010110001;
                8'b11110101 : exp_trans.out_10b = 10'b1010100001;
                8'b11110110 : exp_trans.out_10b = 10'b0110100001;
                8'b11110111 : exp_trans.out_10b = 10'b0001011110;
                8'b11111000 : exp_trans.out_10b = 10'b0011001110;
                8'b11111001 : exp_trans.out_10b = 10'b1001100001;
                8'b11111010 : exp_trans.out_10b = 10'b0101100001;
                8'b11111011 : exp_trans.out_10b = 10'b0010011110;
                8'b11111100 : exp_trans.out_10b = 10'b0011100001;
                8'b11111101 : exp_trans.out_10b = 10'b0100011110;
                8'b11111110 : exp_trans.out_10b = 10'b1000011110;
                8'b11111111 : exp_trans.out_10b = 10'b0101001110;
                default : exp_trans.out_10b = 10'b0000000000;
           endcase
        end
        
        for(int i = 0; i < 10; i++) begin
            rm_queue.push_back(exp_trans.out_10b[i]);
        end
        
        if (exp_trans.out_10b[0]+exp_trans.out_10b[1]+exp_trans.out_10b[2]+exp_trans.out_10b[3]+exp_trans.out_10b[4]+exp_trans.out_10b[5]+exp_trans.out_10b[6]+exp_trans.out_10b[7]+exp_trans.out_10b[8]+exp_trans.out_10b[9] > 5)
          exp_trans.out_RD = 2'sb01; //RD = +1 (more 1s then +1 RD)
        else if (exp_trans.out_10b[0]+exp_trans.out_10b[1]+exp_trans.out_10b[2]+exp_trans.out_10b[3]+exp_trans.out_10b[4]+exp_trans.out_10b[5]+exp_trans.out_10b[6]+exp_trans.out_10b[7]+exp_trans.out_10b[8]+exp_trans.out_10b[9] < 5)
          exp_trans.out_RD = 2'sb11; //RD = -1 (more 0s then -1 RD)
        else
          exp_trans.out_RD = exp_trans.in_RD;
          
        `uvm_info(get_full_name(), $sformatf("EXPECTED TRANSACTION FROM REF MODEL"), UVM_LOW);
        exp_trans.print();
        rm2sb_port.write(exp_trans);
     endtask
endclass

`endif
     
