`ifndef SERDES_REF_MODEL_PKG
`define SERDES_REF_MODEL_PKG

package serdes_ref_model_pkg;
    import uvm_pkg::*;
   `include "uvm_macros.svh"
   
   import serdes_agent_pkg::*;
   
   `include "ser_ref_model.sv"
   
endpackage

`endif
