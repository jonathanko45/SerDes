`ifndef SER_SEQUENCE_LIB
`define SER_SEQUENCE_LIB

package ser_sequence_lib;
   
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import ser_agent_pkg::*;
    import ser_env_pkg::*;
    
    //including ser test list
    `include "ser_random_sequence.sv"
    `include "ser_multiple_random_sequence.sv"
    
endpackage

`endif


